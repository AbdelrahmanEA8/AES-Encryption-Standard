package AES_pack;

    import uvm_pkg::*;
    `include "uvm_macros.svh"
    `include "AES_seq_item.svh"
    `include "AES_sequence.svh"
    `include "AES_driver.svh"
    `include "AES_monitor.svh"
    `include "AES_sequencer.svh"
    `include "AES_agent.svh"
    `include "AES_scoreboard.svh"
    `include "AES_subscriber.svh"
    `include "AES_env.svh"
    `include "AES_test.svh"

endpackage